//------------------------------------------------------------------------------
// Definitions and macros for adder agent
//------------------------------------------------------------------------------
// This file contains definitions and macros used by the adder agent.
//
// Author: Nelson Alves nelsonafn@gmail.com
// Date  : October 2023
//------------------------------------------------------------------------------

`ifndef ADDER_DEFINES
`define ADDER_DEFINES

  `define ADDER_WIDTH 4 
  `define NO_OF_TRANSACTIONS 1000

`endif
